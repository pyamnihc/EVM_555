.title KiCad schematic
.include "D:/hw_things/EVM_555_spice.lib"
.model Q17.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q18.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q16.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q19B1.MMBT3906 PNP
+                     is=6.84896e-14
+                     bf=135.6
+                     nf=1
+                     vaf=18.7
+                     ikf=0.0882
+                     ise=5.52481e-13
+                     ne=1.5
+                     br=0.304
+                     nr=1
+                     var=200
+                     ikr=0.229087
+                     isc=171.764p
+                     nc=1.5
+                     rb=1.05
+                     irb=1.51189m
+                     rbm=0.011
+                     re=0.022
+                     rc=1.57
+                     cje=8.03203p
+                     vje=0.711825
+                     mje=0.304224
+                     tf=319.3p
+                     xtf=6
+                     vtf=4
+                     itf=0.4
+                     cjc=9.50523p
+                     vjc=0.841441
+                     mjc=0.5
+                     tr=33.42n
+                     xtb=1.58
+                     eg=0.78
+                     xti=3
+                     fc=0.5
.model Q9.MMBT3906 PNP
+                  is=6.84896e-14
+                  bf=135.6
+                  nf=1
+                  vaf=18.7
+                  ikf=0.0882
+                  ise=5.52481e-13
+                  ne=1.5
+                  br=0.304
+                  nr=1
+                  var=200
+                  ikr=0.229087
+                  isc=171.764p
+                  nc=1.5
+                  rb=1.05
+                  irb=1.51189m
+                  rbm=0.011
+                  re=0.022
+                  rc=1.57
+                  cje=8.03203p
+                  vje=0.711825
+                  mje=0.304224
+                  tf=319.3p
+                  xtf=6
+                  vtf=4
+                  itf=0.4
+                  cjc=9.50523p
+                  vjc=0.841441
+                  mjc=0.5
+                  tr=33.42n
+                  xtb=1.58
+                  eg=0.78
+                  xti=3
+                  fc=0.5
.model Q10.MMBT3906 PNP
+                   is=6.84896e-14
+                   bf=135.6
+                   nf=1
+                   vaf=18.7
+                   ikf=0.0882
+                   ise=5.52481e-13
+                   ne=1.5
+                   br=0.304
+                   nr=1
+                   var=200
+                   ikr=0.229087
+                   isc=171.764p
+                   nc=1.5
+                   rb=1.05
+                   irb=1.51189m
+                   rbm=0.011
+                   re=0.022
+                   rc=1.57
+                   cje=8.03203p
+                   vje=0.711825
+                   mje=0.304224
+                   tf=319.3p
+                   xtf=6
+                   vtf=4
+                   itf=0.4
+                   cjc=9.50523p
+                   vjc=0.841441
+                   mjc=0.5
+                   tr=33.42n
+                   xtb=1.58
+                   eg=0.78
+                   xti=3
+                   fc=0.5
.model Q20.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q14.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q21.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q19A1.MMBT3906 PNP
+                     is=6.84896e-14
+                     bf=135.6
+                     nf=1
+                     vaf=18.7
+                     ikf=0.0882
+                     ise=5.52481e-13
+                     ne=1.5
+                     br=0.304
+                     nr=1
+                     var=200
+                     ikr=0.229087
+                     isc=171.764p
+                     nc=1.5
+                     rb=1.05
+                     irb=1.51189m
+                     rbm=0.011
+                     re=0.022
+                     rc=1.57
+                     cje=8.03203p
+                     vje=0.711825
+                     mje=0.304224
+                     tf=319.3p
+                     xtf=6
+                     vtf=4
+                     itf=0.4
+                     cjc=9.50523p
+                     vjc=0.841441
+                     mjc=0.5
+                     tr=33.42n
+                     xtb=1.58
+                     eg=0.78
+                     xti=3
+                     fc=0.5
.model Q15.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q11.MMBT3906 PNP
+                   is=6.84896e-14
+                   bf=135.6
+                   nf=1
+                   vaf=18.7
+                   ikf=0.0882
+                   ise=5.52481e-13
+                   ne=1.5
+                   br=0.304
+                   nr=1
+                   var=200
+                   ikr=0.229087
+                   isc=171.764p
+                   nc=1.5
+                   rb=1.05
+                   irb=1.51189m
+                   rbm=0.011
+                   re=0.022
+                   rc=1.57
+                   cje=8.03203p
+                   vje=0.711825
+                   mje=0.304224
+                   tf=319.3p
+                   xtf=6
+                   vtf=4
+                   itf=0.4
+                   cjc=9.50523p
+                   vjc=0.841441
+                   mjc=0.5
+                   tr=33.42n
+                   xtb=1.58
+                   eg=0.78
+                   xti=3
+                   fc=0.5
.model Q13.MMBT3906 PNP
+                   is=6.84896e-14
+                   bf=135.6
+                   nf=1
+                   vaf=18.7
+                   ikf=0.0882
+                   ise=5.52481e-13
+                   ne=1.5
+                   br=0.304
+                   nr=1
+                   var=200
+                   ikr=0.229087
+                   isc=171.764p
+                   nc=1.5
+                   rb=1.05
+                   irb=1.51189m
+                   rbm=0.011
+                   re=0.022
+                   rc=1.57
+                   cje=8.03203p
+                   vje=0.711825
+                   mje=0.304224
+                   tf=319.3p
+                   xtf=6
+                   vtf=4
+                   itf=0.4
+                   cjc=9.50523p
+                   vjc=0.841441
+                   mjc=0.5
+                   tr=33.42n
+                   xtb=1.58
+                   eg=0.78
+                   xti=3
+                   fc=0.5
.model Q12.MMBT3906 PNP
+                   is=6.84896e-14
+                   bf=135.6
+                   nf=1
+                   vaf=18.7
+                   ikf=0.0882
+                   ise=5.52481e-13
+                   ne=1.5
+                   br=0.304
+                   nr=1
+                   var=200
+                   ikr=0.229087
+                   isc=171.764p
+                   nc=1.5
+                   rb=1.05
+                   irb=1.51189m
+                   rbm=0.011
+                   re=0.022
+                   rc=1.57
+                   cje=8.03203p
+                   vje=0.711825
+                   mje=0.304224
+                   tf=319.3p
+                   xtf=6
+                   vtf=4
+                   itf=0.4
+                   cjc=9.50523p
+                   vjc=0.841441
+                   mjc=0.5
+                   tr=33.42n
+                   xtb=1.58
+                   eg=0.78
+                   xti=3
+                   fc=0.5
.model Q19.MMBT3906 PNP
+                   is=6.84896e-14
+                   bf=135.6
+                   nf=1
+                   vaf=18.7
+                   ikf=0.0882
+                   ise=5.52481e-13
+                   ne=1.5
+                   br=0.304
+                   nr=1
+                   var=200
+                   ikr=0.229087
+                   isc=171.764p
+                   nc=1.5
+                   rb=1.05
+                   irb=1.51189m
+                   rbm=0.011
+                   re=0.022
+                   rc=1.57
+                   cje=8.03203p
+                   vje=0.711825
+                   mje=0.304224
+                   tf=319.3p
+                   xtf=6
+                   vtf=4
+                   itf=0.4
+                   cjc=9.50523p
+                   vjc=0.841441
+                   mjc=0.5
+                   tr=33.42n
+                   xtb=1.58
+                   eg=0.78
+                   xti=3
+                   fc=0.5
.model Q22.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q24.MMBT3904 NPN
+                   is=4.639e-15
+                   bf=160.1
+                   nf=0.9995
+                   vaf=98.69
+                   ikf=0.12
+                   ise=2.091e-14
+                   ne=1.6
+                   br=5.944
+                   nr=1.001
+                   var=19.29
+                   ikr=0.06
+                   isc=3.257p
+                   nc=1.394
+                   rb=1
+                   re=0.3614
+                   rc=1.755
+                   cje=5.631p
+                   vje=0.7002
+                   mje=0.3385
+                   tf=300.1p
+                   xtf=27
+                   vtf=1.461
+                   itf=0.2723
+                   cjc=4.949p
+                   vjc=0.5969
+                   mjc=0.1928
+                   xcjc=0.864
+                   tr=94n
+                   xtb=0
+                   eg=1.11
+                   xti=3
+                   fc=0.5582
.model Q23.MMBT3906 PNP
+                   is=6.84896e-14
+                   bf=135.6
+                   nf=1
+                   vaf=18.7
+                   ikf=0.0882
+                   ise=5.52481e-13
+                   ne=1.5
+                   br=0.304
+                   nr=1
+                   var=200
+                   ikr=0.229087
+                   isc=171.764p
+                   nc=1.5
+                   rb=1.05
+                   irb=1.51189m
+                   rbm=0.011
+                   re=0.022
+                   rc=1.57
+                   cje=8.03203p
+                   vje=0.711825
+                   mje=0.304224
+                   tf=319.3p
+                   xtf=6
+                   vtf=4
+                   itf=0.4
+                   cjc=9.50523p
+                   vjc=0.841441
+                   mjc=0.5
+                   tr=33.42n
+                   xtb=1.58
+                   eg=0.78
+                   xti=3
+                   fc=0.5
.model Q4.MMBT3904 NPN
+                  is=4.639e-15
+                  bf=160.1
+                  nf=0.9995
+                  vaf=98.69
+                  ikf=0.12
+                  ise=2.091e-14
+                  ne=1.6
+                  br=5.944
+                  nr=1.001
+                  var=19.29
+                  ikr=0.06
+                  isc=3.257p
+                  nc=1.394
+                  rb=1
+                  re=0.3614
+                  rc=1.755
+                  cje=5.631p
+                  vje=0.7002
+                  mje=0.3385
+                  tf=300.1p
+                  xtf=27
+                  vtf=1.461
+                  itf=0.2723
+                  cjc=4.949p
+                  vjc=0.5969
+                  mjc=0.1928
+                  xcjc=0.864
+                  tr=94n
+                  xtb=0
+                  eg=1.11
+                  xti=3
+                  fc=0.5582
.model Q3.MMBT3904 NPN
+                  is=4.639e-15
+                  bf=160.1
+                  nf=0.9995
+                  vaf=98.69
+                  ikf=0.12
+                  ise=2.091e-14
+                  ne=1.6
+                  br=5.944
+                  nr=1.001
+                  var=19.29
+                  ikr=0.06
+                  isc=3.257p
+                  nc=1.394
+                  rb=1
+                  re=0.3614
+                  rc=1.755
+                  cje=5.631p
+                  vje=0.7002
+                  mje=0.3385
+                  tf=300.1p
+                  xtf=27
+                  vtf=1.461
+                  itf=0.2723
+                  cjc=4.949p
+                  vjc=0.5969
+                  mjc=0.1928
+                  xcjc=0.864
+                  tr=94n
+                  xtb=0
+                  eg=1.11
+                  xti=3
+                  fc=0.5582
.model Q7.MMBT3906 PNP
+                  is=6.84896e-14
+                  bf=135.6
+                  nf=1
+                  vaf=18.7
+                  ikf=0.0882
+                  ise=5.52481e-13
+                  ne=1.5
+                  br=0.304
+                  nr=1
+                  var=200
+                  ikr=0.229087
+                  isc=171.764p
+                  nc=1.5
+                  rb=1.05
+                  irb=1.51189m
+                  rbm=0.011
+                  re=0.022
+                  rc=1.57
+                  cje=8.03203p
+                  vje=0.711825
+                  mje=0.304224
+                  tf=319.3p
+                  xtf=6
+                  vtf=4
+                  itf=0.4
+                  cjc=9.50523p
+                  vjc=0.841441
+                  mjc=0.5
+                  tr=33.42n
+                  xtb=1.58
+                  eg=0.78
+                  xti=3
+                  fc=0.5
.model Q1.MMBT3904 NPN
+                  is=4.639e-15
+                  bf=160.1
+                  nf=0.9995
+                  vaf=98.69
+                  ikf=0.12
+                  ise=2.091e-14
+                  ne=1.6
+                  br=5.944
+                  nr=1.001
+                  var=19.29
+                  ikr=0.06
+                  isc=3.257p
+                  nc=1.394
+                  rb=1
+                  re=0.3614
+                  rc=1.755
+                  cje=5.631p
+                  vje=0.7002
+                  mje=0.3385
+                  tf=300.1p
+                  xtf=27
+                  vtf=1.461
+                  itf=0.2723
+                  cjc=4.949p
+                  vjc=0.5969
+                  mjc=0.1928
+                  xcjc=0.864
+                  tr=94n
+                  xtb=0
+                  eg=1.11
+                  xti=3
+                  fc=0.5582
.model Q6.MMBT3906 PNP
+                  is=6.84896e-14
+                  bf=135.6
+                  nf=1
+                  vaf=18.7
+                  ikf=0.0882
+                  ise=5.52481e-13
+                  ne=1.5
+                  br=0.304
+                  nr=1
+                  var=200
+                  ikr=0.229087
+                  isc=171.764p
+                  nc=1.5
+                  rb=1.05
+                  irb=1.51189m
+                  rbm=0.011
+                  re=0.022
+                  rc=1.57
+                  cje=8.03203p
+                  vje=0.711825
+                  mje=0.304224
+                  tf=319.3p
+                  xtf=6
+                  vtf=4
+                  itf=0.4
+                  cjc=9.50523p
+                  vjc=0.841441
+                  mjc=0.5
+                  tr=33.42n
+                  xtb=1.58
+                  eg=0.78
+                  xti=3
+                  fc=0.5
.model Q5.MMBT3906 PNP
+                  is=6.84896e-14
+                  bf=135.6
+                  nf=1
+                  vaf=18.7
+                  ikf=0.0882
+                  ise=5.52481e-13
+                  ne=1.5
+                  br=0.304
+                  nr=1
+                  var=200
+                  ikr=0.229087
+                  isc=171.764p
+                  nc=1.5
+                  rb=1.05
+                  irb=1.51189m
+                  rbm=0.011
+                  re=0.022
+                  rc=1.57
+                  cje=8.03203p
+                  vje=0.711825
+                  mje=0.304224
+                  tf=319.3p
+                  xtf=6
+                  vtf=4
+                  itf=0.4
+                  cjc=9.50523p
+                  vjc=0.841441
+                  mjc=0.5
+                  tr=33.42n
+                  xtb=1.58
+                  eg=0.78
+                  xti=3
+                  fc=0.5
.model Q8.MMBT3906 PNP
+                  is=6.84896e-14
+                  bf=135.6
+                  nf=1
+                  vaf=18.7
+                  ikf=0.0882
+                  ise=5.52481e-13
+                  ne=1.5
+                  br=0.304
+                  nr=1
+                  var=200
+                  ikr=0.229087
+                  isc=171.764p
+                  nc=1.5
+                  rb=1.05
+                  irb=1.51189m
+                  rbm=0.011
+                  re=0.022
+                  rc=1.57
+                  cje=8.03203p
+                  vje=0.711825
+                  mje=0.304224
+                  tf=319.3p
+                  xtf=6
+                  vtf=4
+                  itf=0.4
+                  cjc=9.50523p
+                  vjc=0.841441
+                  mjc=0.5
+                  tr=33.42n
+                  xtb=1.58
+                  eg=0.78
+                  xti=3
+                  fc=0.5
.model Q2.MMBT3904 NPN
+                  is=4.639e-15
+                  bf=160.1
+                  nf=0.9995
+                  vaf=98.69
+                  ikf=0.12
+                  ise=2.091e-14
+                  ne=1.6
+                  br=5.944
+                  nr=1.001
+                  var=19.29
+                  ikr=0.06
+                  isc=3.257p
+                  nc=1.394
+                  rb=1
+                  re=0.3614
+                  rc=1.755
+                  cje=5.631p
+                  vje=0.7002
+                  mje=0.3385
+                  tf=300.1p
+                  xtf=27
+                  vtf=1.461
+                  itf=0.2723
+                  cjc=4.949p
+                  vjc=0.5969
+                  mjc=0.1928
+                  xcjc=0.864
+                  tr=94n
+                  xtb=0
+                  eg=1.11
+                  xti=3
+                  fc=0.5582
.save all
.probe alli
R16 Net-_Q20-E_ Net-_Q19-C_ 100
R15 Net-_Q20-E_ GND 4.7k
R11 Net-_Q17-C_ thresh_out 4.7k
Q17 Net-_Q16-C_ GND Net-_Q17-C_ Q17.MMBT3904
Q18 Net-_Q18-B_ Net-_Q16-C_ Net-_Q18-B_ Q18.MMBT3904
Q16 thresh_out GND Net-_Q16-C_ Q16.MMBT3904
R10 Net-_Q19A1-B_ Net-_Q18-B_ 15k
Q19B1 Net-_Q19A1-B_ VCC Net-_Q19A1-B_ Q19B1.MMBT3906
Q9 Net-_Q19A1-B_ Net-_Q9-E_ Net-_Q10-E_ Q9.MMBT3906
Q10 Net-_Q10-B_ Net-_Q10-E_ GND Q10.MMBT3906
R4 VCC Net-_Q9-E_ 1k
Q20 Net-_Q17-C_ Net-_Q20-E_ Net-_Q20-C_ Q20.MMBT3904
R12 VCC Net-_Q20-C_ 6.8k
R13 Net-_Q14-B_ Net-_J11-Pin_1_ 3.9k
Q14 Net-_Q14-B_ Net-_J11-Pin_1_ VCC Q14.MMBT3904
Q21 Net-_Q20-C_ Net-_Q14-B_ VCC Q21.MMBT3904
Q19A1 Net-_Q19A1-B_ VCC Net-_Q17-C_ Q19A1.MMBT3906
R6 Net-_Q12-C_ GND 100k
Q15 Net-_Q12-C_ GND thresh_out Q15.MMBT3904
Q11 Net-_Q11-B_ Net-_Q10-B_ GND Q11.MMBT3906
Q13 Net-_J10-Pin_1_ Net-_Q12-B_ GND Q13.MMBT3906
Q12 Net-_Q12-B_ Net-_Q10-E_ Net-_Q12-C_ Q12.MMBT3906
Q19 Net-_Q19-B_ Net-_Q18-B_ Net-_Q19-C_ Q19.MMBT3906
Q22 Net-_Q19-C_ GND Net-_J15-Pin_1_ Q22.MMBT3904
R17 Net-_Q19-B_ Net-_J13-Pin_1_ 100k
Q24 Net-_Q24-B_ GND Net-_J11-Pin_1_ Q24.MMBT3904
Q23 Net-_Q20-C_ Net-_J11-Pin_1_ Net-_Q20-C_ Q23.MMBT3906
R14 Net-_Q20-E_ Net-_Q24-B_ 220
R2 VCC Net-_Q5-E_ 820
Q4 Net-_J7-Pin_1_ Net-_Q3-B_ Net-_Q3-C_ Q4.MMBT3904
Q3 Net-_Q3-B_ Net-_Q2-E_ Net-_Q3-C_ Q3.MMBT3904
Q7 Net-_Q3-C_ Net-_Q5-E_ GND Q7.MMBT3906
Q1 Net-_J5-Pin_1_ Net-_Q1-E_ Net-_Q1-C_ Q1.MMBT3904
Q6 Net-_Q1-C_ Net-_Q6-E_ Net-_Q1-C_ Q6.MMBT3906
Q5 Net-_Q1-C_ Net-_Q5-E_ thresh_out Q5.MMBT3906
R1 VCC Net-_Q6-E_ 4.7k
Q8 Net-_Q3-C_ Net-_Q8-E_ Net-_Q3-C_ Q8.MMBT3906
R8 Net-_J7-Pin_1_ Net-_Q11-B_ 4.7k
R7 VCC Net-_J7-Pin_1_ 4.7k
R3 VCC Net-_Q8-E_ 4.7k
Q2 Net-_Q1-E_ Net-_Q2-E_ Net-_Q1-C_ Q2.MMBT3904
J4 __J4
J3 __J3
R5 Net-_Q2-E_ GND 10k
V1 VCC GND DC 12 
R9 Net-_Q11-B_ GND 4.7k
.end
